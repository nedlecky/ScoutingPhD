module alu4 ( 
	a,
	b,
	sel,
	cin,
	c,
	cout,
	z
	) ;

inout [3:0] a;
inout [3:0] b;
inout [3:0] sel;
inout  cin;
inout [3:0] c;
inout  cout;
inout  z;
res��@ K