LIBRARY IEEE;
USE  IEEE.STD_LOGIC_1164.all;
ENTITY andgate IS
	PORT(
		PB1, PB2		: IN	STD_LOGIC;
		LED				: OUT	STD_LOGIC);
END andgate;
ARCHITECTURE a OF andgate IS
BEGIN
	LED <= PB1 AND PB2;
END a;

