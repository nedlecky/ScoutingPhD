-- 5-bit x 5-bit Signed Multiplier
-- Direct TT Implementation of [B&V] algorithm

-- University of Vermont
-- EE 231: Digital Computer Design I Spring 2002
-- Dr. Ned Lecky

library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_arith.all;
use ieee.std_logic_unsigned.all;

entity multiplier is
	port
	(
		x_in,y_in	: in	std_logic_vector(4 downto 0);
		f			: out	std_logic_vector(9 downto 0)
	);
end multiplier;

architecture arch of multiplier is
	signal inputs : integer range 0 to 1023;
begin
	inputs <= conv_integer(x_in & y_in);
        with inputs select
        f(0) <= '1' when
        33|35|37|39|41|43|45|47|49|51|53|55|57|59|61|63|97|99|101|103|105
        |107|109|111|113|115|117|119|121|123|125|127|161|163|165|167|169|171|173|175|177|179
        |181|183|185|187|189|191|225|227|229|231|233|235|237|239|241|243|245|247|249|251|253
        |255|289|291|293|295|297|299|301|303|305|307|309|311|313|315|317|319|353|355|357|359
        |361|363|365|367|369|371|373|375|377|379|381|383|417|419|421|423|425|427|429|431|433
        |435|437|439|441|443|445|447|481|483|485|487|489|491|493|495|497|499|501|503|505|507
        |509|511|545|547|549|551|553|555|557|559|561|563|565|567|569|571|573|575|609|611|613
        |615|617|619|621|623|625|627|629|631|633|635|637|639|673|675|677|679|681|683|685|687
        |689|691|693|695|697|699|701|703|737|739|741|743|745|747|749|751|753|755|757|759|761
        |763|765|767|801|803|805|807|809|811|813|815|817|819|821|823|825|827|829|831|865|867
        |869|871|873|875|877|879|881|883|885|887|889|891|893|895|929|931|933|935|937|939|941
        |943|945|947|949|951|953|955|957|959|993|995|997|999|1001|1003|1005|1007|1009|1011|1013|1015
        |1017|1019|1021|1023,
        '0' when others;

        with inputs select
        f(1) <= '1' when
        34|35|38|39|42|43|46|47|50|51|54|55|58|59|62|63|65|67|69|71|73
        |75|77|79|81|83|85|87|89|91|93|95|97|98|101|102|105|106|109|110|113|114
        |117|118|121|122|125|126|162|163|166|167|170|171|174|175|178|179|182|183|186|187|190
        |191|193|195|197|199|201|203|205|207|209|211|213|215|217|219|221|223|225|226|229|230
        |233|234|237|238|241|242|245|246|249|250|253|254|290|291|294|295|298|299|302|303|306
        |307|310|311|314|315|318|319|321|323|325|327|329|331|333|335|337|339|341|343|345|347
        |349|351|353|354|357|358|361|362|365|366|369|370|373|374|377|378|381|382|418|419|422
        |423|426|427|430|431|434|435|438|439|442|443|446|447|449|451|453|455|457|459|461|463
        |465|467|469|471|473|475|477|479|481|482|485|486|489|490|493|494|497|498|501|502|505
        |506|509|510|546|547|550|551|554|555|558|559|562|563|566|567|570|571|574|575|577|579
        |581|583|585|587|589|591|593|595|597|599|601|603|605|607|609|610|613|614|617|618|621
        |622|625|626|629|630|633|634|637|638|674|675|678|679|682|683|686|687|690|691|694|695
        |698|699|702|703|705|707|709|711|713|715|717|719|721|723|725|727|729|731|733|735|737
        |738|741|742|745|746|749|750|753|754|757|758|761|762|765|766|802|803|806|807|810|811
        |814|815|818|819|822|823|826|827|830|831|833|835|837|839|841|843|845|847|849|851|853
        |855|857|859|861|863|865|866|869|870|873|874|877|878|881|882|885|886|889|890|893|894
        |930|931|934|935|938|939|942|943|946|947|950|951|954|955|958|959|961|963|965|967|969
        |971|973|975|977|979|981|983|985|987|989|991|993|994|997|998|1001|1002|1005|1006|1009|1010
        |1013|1014|1017|1018|1021|1022,
        '0' when others;

        with inputs select
        f(2) <= '1' when
        36|37|38|39|44|45|46|47|52|53|54|55|60|61|62|63|66|67|70|71|74
        |75|78|79|82|83|86|87|90|91|94|95|98|100|101|103|106|108|109|111|114|116
        |117|119|122|124|125|127|129|131|133|135|137|139|141|143|145|147|149|151|153|155|157
        |159|161|163|164|166|169|171|172|174|177|179|180|182|185|187|188|190|193|194|197|198
        |201|202|205|206|209|210|213|214|217|218|221|222|225|226|227|228|233|234|235|236|241
        |242|243|244|249|250|251|252|292|293|294|295|300|301|302|303|308|309|310|311|316|317
        |318|319|322|323|326|327|330|331|334|335|338|339|342|343|346|347|350|351|354|356|357
        |359|362|364|365|367|370|372|373|375|378|380|381|383|385|387|389|391|393|395|397|399
        |401|403|405|407|409|411|413|415|417|419|420|422|425|427|428|430|433|435|436|438|441
        |443|444|446|449|450|453|454|457|458|461|462|465|466|469|470|473|474|477|478|481|482
        |483|484|489|490|491|492|497|498|499|500|505|506|507|508|548|549|550|551|556|557|558
        |559|564|565|566|567|572|573|574|575|578|579|582|583|586|587|590|591|594|595|598|599
        |602|603|606|607|610|612|613|615|618|620|621|623|626|628|629|631|634|636|637|639|641
        |643|645|647|649|651|653|655|657|659|661|663|665|667|669|671|673|675|676|678|681|683
        |684|686|689|691|692|694|697|699|700|702|705|706|709|710|713|714|717|718|721|722|725
        |726|729|730|733|734|737|738|739|740|745|746|747|748|753|754|755|756|761|762|763|764
        |804|805|806|807|812|813|814|815|820|821|822|823|828|829|830|831|834|835|838|839|842
        |843|846|847|850|851|854|855|858|859|862|863|866|868|869|871|874|876|877|879|882|884
        |885|887|890|892|893|895|897|899|901|903|905|907|909|911|913|915|917|919|921|923|925
        |927|929|931|932|934|937|939|940|942|945|947|948|950|953|955|956|958|961|962|965|966
        |969|970|973|974|977|978|981|982|985|986|989|990|993|994|995|996|1001|1002|1003|1004|1009
        |1010|1011|1012|1017|1018|1019|1020,
        '0' when others;

        with inputs select
        f(3) <= '1' when
        40|41|42|43|44|45|46|47|56|57|58|59|60|61|62|63|68|69|70|71|76
        |77|78|79|84|85|86|87|92|93|94|95|99|100|101|104|105|106|110|111|115|116
        |117|120|121|122|126|127|130|131|134|135|138|139|142|143|146|147|150|151|154|155|158
        |159|162|163|165|166|168|169|172|175|178|179|181|182|184|185|188|191|194|196|197|199
        |202|204|205|207|210|212|213|215|218|220|221|223|226|228|230|232|233|235|237|239|242
        |244|246|248|249|251|253|255|257|259|261|263|265|267|269|271|273|275|277|279|281|283
        |285|287|289|291|293|295|296|298|300|302|305|307|309|311|312|314|316|318|321|323|324
        |326|329|331|332|334|337|339|340|342|345|347|348|350|353|356|359|360|362|363|365|366
        |369|372|375|376|378|379|381|382|385|386|389|390|393|394|397|398|401|402|405|406|409
        |410|413|414|417|418|422|423|424|427|428|429|433|434|438|439|440|443|444|445|449|450
        |451|452|457|458|459|460|465|466|467|468|473|474|475|476|481|482|483|484|485|486|487
        |488|497|498|499|500|501|502|503|504|552|553|554|555|556|557|558|559|568|569|570|571
        |572|573|574|575|580|581|582|583|588|589|590|591|596|597|598|599|604|605|606|607|611
        |612|613|616|617|618|622|623|627|628|629|632|633|634|638|639|642|643|646|647|650|651
        |654|655|658|659|662|663|666|667|670|671|674|675|677|678|680|681|684|687|690|691|693
        |694|696|697|700|703|706|708|709|711|714|716|717|719|722|724|725|727|730|732|733|735
        |738|740|742|744|745|747|749|751|754|756|758|760|761|763|765|767|769|771|773|775|777
        |779|781|783|785|787|789|791|793|795|797|799|801|803|805|807|808|810|812|814|817|819
        |821|823|824|826|828|830|833|835|836|838|841|843|844|846|849|851|852|854|857|859|860
        |862|865|868|871|872|874|875|877|878|881|884|887|888|890|891|893|894|897|898|901|902
        |905|906|909|910|913|914|917|918|921|922|925|926|929|930|934|935|936|939|940|941|945
        |946|950|951|952|955|956|957|961|962|963|964|969|970|971|972|977|978|979|980|985|986
        |987|988|993|994|995|996|997|998|999|1000|1009|1010|1011|1012|1013|1014|1015|1016,
        '0' when others;

        with inputs select
        f(4) <= '1' when
        48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|72|73|74|75|76
        |77|78|79|88|89|90|91|92|93|94|95|102|103|104|105|106|112|113|114|115|116
        |117|123|124|125|126|127|132|133|134|135|140|141|142|143|148|149|150|151|156|157|158
        |159|164|165|166|170|171|172|176|177|178|179|183|184|185|189|190|191|195|196|197|200
        |201|202|206|207|211|212|213|216|217|218|222|223|227|228|231|232|233|236|237|240|241
        |242|245|246|250|251|254|255|258|259|262|263|266|267|270|271|274|275|278|279|282|283
        |286|287|290|291|294|295|297|298|301|302|304|305|308|309|312|315|316|319|322|323|325
        |326|328|329|332|335|338|339|341|342|344|345|348|351|354|357|360|363|366|368|369|371
        |372|374|375|377|378|380|381|383|386|388|389|391|394|396|397|399|402|404|405|407|410
        |412|413|415|418|420|423|425|428|430|432|433|435|437|438|440|442|443|445|447|450|452
        |454|456|457|459|461|463|466|468|470|472|473|475|477|479|482|484|486|488|490|492|494
        |496|497|499|501|503|505|507|509|511|513|515|517|519|521|523|525|527|529|531|533|535
        |537|539|541|543|545|547|549|551|553|555|557|559|560|562|564|566|568|570|572|574|577
        |579|581|583|584|586|588|590|593|595|597|599|600|602|604|606|609|611|613|614|616|618
        |619|621|623|624|626|628|631|633|636|638|641|643|644|646|649|651|652|654|657|659|660
        |662|665|667|668|670|673|675|676|678|679|681|682|684|685|687|688|690|693|696|699|702
        |705|708|711|712|714|715|717|718|721|724|727|728|730|731|733|734|737|740|741|744|747
        |748|751|752|754|755|758|759|761|762|765|766|769|770|773|774|777|778|781|782|785|786
        |789|790|793|794|797|798|801|802|805|806|810|811|814|815|816|819|820|823|824|825|828
        |829|833|834|838|839|840|843|844|845|849|850|854|855|856|859|860|861|865|866|867|871
        |872|873|877|878|879|880|884|885|886|890|891|892|897|898|899|900|905|906|907|908|913
        |914|915|916|921|922|923|924|929|930|931|932|933|939|940|941|942|943|944|950|951|952
        |953|954|961|962|963|964|965|966|967|968|977|978|979|980|981|982|983|984|993|994|995
        |996|997|998|999|1000|1001|1002|1003|1004|1005|1006|1007|1008,
        '0' when others;

        with inputs select
        f(5) <= '1' when
        48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|80|81|82|83|84
        |85|86|87|88|89|90|91|92|93|94|95|107|108|109|110|111|118|119|120|121|122
        |123|124|125|126|127|136|137|138|139|140|141|142|143|152|153|154|155|156|157|158|159
        |167|168|169|170|171|172|176|177|178|179|186|187|188|189|190|191|198|199|200|201|202
        |208|209|210|211|212|213|219|220|221|222|223|229|230|231|232|233|238|239|243|244|245
        |246|252|253|254|255|260|261|262|263|268|269|270|271|276|277|278|279|284|285|286|287
        |292|293|294|295|299|300|301|302|304|305|310|311|312|317|318|319|324|325|326|330|331
        |332|336|337|338|339|343|344|345|349|350|351|355|356|357|361|362|363|367|370|371|372
        |376|377|378|382|383|387|388|389|392|393|394|398|399|403|404|405|408|409|410|414|415
        |419|420|424|425|429|430|432|433|436|437|438|441|442|443|446|447|451|452|455|456|457
        |460|461|464|465|466|469|470|474|475|478|479|483|484|487|488|491|492|495|498|499|502
        |503|506|507|510|511|513|514|517|518|521|522|525|526|529|530|533|534|537|538|541|542
        |545|546|549|550|553|554|557|558|560|561|564|565|568|569|572|573|577|578|581|582|586
        |587|590|591|592|595|596|599|600|601|604|605|609|610|613|614|615|618|619|620|623|626
        |627|631|632|636|637|641|642|646|647|648|651|652|653|657|658|662|663|664|667|668|669
        |673|674|678|679|680|684|685|686|688|689|693|694|695|699|700|701|705|706|707|711|712
        |713|717|718|719|720|724|725|726|730|731|732|737|738|739|744|745|746|751|754|755|756
        |757|761|762|763|764|769|770|771|772|777|778|779|780|785|786|787|788|793|794|795|796
        |801|802|803|804|810|811|812|813|816|817|818|823|824|825|826|827|833|834|835|836|837
        |843|844|845|846|847|848|854|855|856|857|858|865|866|867|868|869|870|877|878|879|884
        |885|886|887|888|889|897|898|899|900|901|902|903|904|913|914|915|916|917|918|919|920
        |929|930|931|932|933|934|935|936|937|938|944|945|946|947|948|949|961|962|963|964|965
        |966|967|968|969|970|971|972|973|974|975|976|993|994|995|996|997|998|999|1000|1001|1002
        |1003|1004|1005|1006|1007,
        '0' when others;

        with inputs select
        f(6) <= '1' when
        48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|80|81|82|83|84
        |85|86|87|88|89|90|91|92|93|94|95|112|113|114|115|116|117|118|119|120|121
        |122|123|124|125|126|127|144|145|146|147|148|149|150|151|152|153|154|155|156|157|158
        |159|173|174|175|180|181|182|183|184|185|186|187|188|189|190|191|203|204|205|206|207
        |214|215|216|217|218|219|220|221|222|223|234|235|236|237|238|239|247|248|249|250|251
        |252|253|254|255|264|265|266|267|268|269|270|271|280|281|282|283|284|285|286|287|296
        |297|298|299|300|301|302|304|305|313|314|315|316|317|318|319|327|328|329|330|331|332
        |336|337|338|339|346|347|348|349|350|351|358|359|360|361|362|363|368|369|370|371|372
        |379|380|381|382|383|390|391|392|393|394|400|401|402|403|404|405|411|412|413|414|415
        |421|422|423|424|425|431|434|435|436|437|438|444|445|446|447|453|454|455|456|457|462
        |463|467|468|469|470|476|477|478|479|485|486|487|488|493|494|495|500|501|502|503|508
        |509|510|511|513|514|515|516|521|522|523|524|529|530|531|532|537|538|539|540|545|546
        |547|548|553|554|555|556|560|561|562|563|568|569|570|571|577|578|579|580|586|587|588
        |589|592|593|594|599|600|601|602|603|609|610|611|612|618|619|620|621|622|624|625|631
        |632|633|634|635|641|642|643|644|645|651|652|653|654|655|656|662|663|664|665|666|673
        |674|675|676|677|684|685|686|687|693|694|695|696|697|698|705|706|707|708|709|710|717
        |718|719|724|725|726|727|728|729|737|738|739|740|741|742|743|751|754|755|756|757|758
        |759|760|769|770|771|772|773|774|775|776|785|786|787|788|789|790|791|792|801|802|803
        |804|805|806|807|808|809|816|817|818|819|820|821|822|833|834|835|836|837|838|839|840
        |841|842|848|849|850|851|852|853|865|866|867|868|869|870|871|872|873|874|875|876|880
        |881|882|883|897|898|899|900|901|902|903|904|905|906|907|908|909|910|911|912|929|930
        |931|932|933|934|935|936|937|938|939|940|941|942|943|961|962|963|964|965|966|967|968
        |969|970|971|972|973|974|975|993|994|995|996|997|998|999|1000|1001|1002|1003|1004|1005|1006
        |1007,
        '0' when others;

        with inputs select
        f(7) <= '1' when
        48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|80|81|82|83|84
        |85|86|87|88|89|90|91|92|93|94|95|112|113|114|115|116|117|118|119|120|121
        |122|123|124|125|126|127|144|145|146|147|148|149|150|151|152|153|154|155|156|157|158
        |159|176|177|178|179|180|181|182|183|184|185|186|187|188|189|190|191|208|209|210|211
        |212|213|214|215|216|217|218|219|220|221|222|223|240|241|242|243|244|245|246|247|248
        |249|250|251|252|253|254|255|272|273|274|275|276|277|278|279|280|281|282|283|284|285
        |286|287|303|306|307|308|309|310|311|312|313|314|315|316|317|318|319|333|334|335|340
        |341|342|343|344|345|346|347|348|349|350|351|364|365|366|367|373|374|375|376|377|378
        |379|380|381|382|383|395|396|397|398|399|406|407|408|409|410|411|412|413|414|415|426
        |427|428|429|430|431|439|440|441|442|443|444|445|446|447|458|459|460|461|462|463|471
        |472|473|474|475|476|477|478|479|489|490|491|492|493|494|495|504|505|506|507|508|509
        |510|511|513|514|515|516|517|518|519|520|529|530|531|532|533|534|535|536|545|546|547
        |548|549|550|551|552|560|561|562|563|564|565|566|567|577|578|579|580|581|582|583|584
        |585|592|593|594|595|596|597|598|609|610|611|612|613|614|615|616|617|624|625|626|627
        |628|629|630|641|642|643|644|645|646|647|648|649|650|656|657|658|659|660|661|673|674
        |675|676|677|678|679|680|681|682|683|688|689|690|691|692|705|706|707|708|709|710|711
        |712|713|714|715|716|720|721|722|723|737|738|739|740|741|742|743|744|745|746|747|748
        |749|750|752|753|769|770|771|772|773|774|775|776|777|778|779|780|781|782|783|784|801
        |802|803|804|805|806|807|808|809|810|811|812|813|814|815|833|834|835|836|837|838|839
        |840|841|842|843|844|845|846|847|865|866|867|868|869|870|871|872|873|874|875|876|877
        |878|879|897|898|899|900|901|902|903|904|905|906|907|908|909|910|911|929|930|931|932
        |933|934|935|936|937|938|939|940|941|942|943|961|962|963|964|965|966|967|968|969|970
        |971|972|973|974|975|993|994|995|996|997|998|999|1000|1001|1002|1003|1004|1005|1006|1007,
        '0' when others;

        with inputs select
        f(8) <= '1' when
        48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|80|81|82|83|84
        |85|86|87|88|89|90|91|92|93|94|95|112|113|114|115|116|117|118|119|120|121
        |122|123|124|125|126|127|144|145|146|147|148|149|150|151|152|153|154|155|156|157|158
        |159|176|177|178|179|180|181|182|183|184|185|186|187|188|189|190|191|208|209|210|211
        |212|213|214|215|216|217|218|219|220|221|222|223|240|241|242|243|244|245|246|247|248
        |249|250|251|252|253|254|255|272|273|274|275|276|277|278|279|280|281|282|283|284|285
        |286|287|304|305|306|307|308|309|310|311|312|313|314|315|316|317|318|319|336|337|338
        |339|340|341|342|343|344|345|346|347|348|349|350|351|368|369|370|371|372|373|374|375
        |376|377|378|379|380|381|382|383|400|401|402|403|404|405|406|407|408|409|410|411|412
        |413|414|415|432|433|434|435|436|437|438|439|440|441|442|443|444|445|446|447|464|465
        |466|467|468|469|470|471|472|473|474|475|476|477|478|479|496|497|498|499|500|501|502
        |503|504|505|506|507|508|509|510|511|513|514|515|516|517|518|519|520|521|522|523|524
        |525|526|527|528|545|546|547|548|549|550|551|552|553|554|555|556|557|558|559|577|578
        |579|580|581|582|583|584|585|586|587|588|589|590|591|609|610|611|612|613|614|615|616
        |617|618|619|620|621|622|623|641|642|643|644|645|646|647|648|649|650|651|652|653|654
        |655|673|674|675|676|677|678|679|680|681|682|683|684|685|686|687|705|706|707|708|709
        |710|711|712|713|714|715|716|717|718|719|737|738|739|740|741|742|743|744|745|746|747
        |748|749|750|751|769|770|771|772|773|774|775|776|777|778|779|780|781|782|783|801|802
        |803|804|805|806|807|808|809|810|811|812|813|814|815|833|834|835|836|837|838|839|840
        |841|842|843|844|845|846|847|865|866|867|868|869|870|871|872|873|874|875|876|877|878
        |879|897|898|899|900|901|902|903|904|905|906|907|908|909|910|911|929|930|931|932|933
        |934|935|936|937|938|939|940|941|942|943|961|962|963|964|965|966|967|968|969|970|971
        |972|973|974|975|993|994|995|996|997|998|999|1000|1001|1002|1003|1004|1005|1006|1007,
        '0' when others;

        with inputs select
        f(9) <= '1' when
        48|49|50|51|52|53|54|55|56|57|58|59|60|61|62|63|80|81|82|83|84
        |85|86|87|88|89|90|91|92|93|94|95|112|113|114|115|116|117|118|119|120|121
        |122|123|124|125|126|127|144|145|146|147|148|149|150|151|152|153|154|155|156|157|158
        |159|176|177|178|179|180|181|182|183|184|185|186|187|188|189|190|191|208|209|210|211
        |212|213|214|215|216|217|218|219|220|221|222|223|240|241|242|243|244|245|246|247|248
        |249|250|251|252|253|254|255|272|273|274|275|276|277|278|279|280|281|282|283|284|285
        |286|287|304|305|306|307|308|309|310|311|312|313|314|315|316|317|318|319|336|337|338
        |339|340|341|342|343|344|345|346|347|348|349|350|351|368|369|370|371|372|373|374|375
        |376|377|378|379|380|381|382|383|400|401|402|403|404|405|406|407|408|409|410|411|412
        |413|414|415|432|433|434|435|436|437|438|439|440|441|442|443|444|445|446|447|464|465
        |466|467|468|469|470|471|472|473|474|475|476|477|478|479|496|497|498|499|500|501|502
        |503|504|505|506|507|508|509|510|511|513|514|515|516|517|518|519|520|521|522|523|524
        |525|526|527|545|546|547|548|549|550|551|552|553|554|555|556|557|558|559|577|578|579
        |580|581|582|583|584|585|586|587|588|589|590|591|609|610|611|612|613|614|615|616|617
        |618|619|620|621|622|623|641|642|643|644|645|646|647|648|649|650|651|652|653|654|655
        |673|674|675|676|677|678|679|680|681|682|683|684|685|686|687|705|706|707|708|709|710
        |711|712|713|714|715|716|717|718|719|737|738|739|740|741|742|743|744|745|746|747|748
        |749|750|751|769|770|771|772|773|774|775|776|777|778|779|780|781|782|783|801|802|803
        |804|805|806|807|808|809|810|811|812|813|814|815|833|834|835|836|837|838|839|840|841
        |842|843|844|845|846|847|865|866|867|868|869|870|871|872|873|874|875|876|877|878|879
        |897|898|899|900|901|902|903|904|905|906|907|908|909|910|911|929|930|931|932|933|934
        |935|936|937|938|939|940|941|942|943|961|962|963|964|965|966|967|968|969|970|971|972
        |973|974|975|993|994|995|996|997|998|999|1000|1001|1002|1003|1004|1005|1006|1007,
        '0' when others;
end arch;

