LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.all;

ENTITY orgate IS
	PORT(
		PB1, PB2	: IN	STD_LOGIC;
		LED		 	: OUT	STD_LOGIC );
END orgate;

ARCHITECTURE a OF orgate IS
BEGIN
	LED <= NOT( NOT PB1 OR NOT PB2 )
END a;


